//: version "1.8.7"

module full_adder(Cout, Cin, B, S, A);
//: interface  /sz:(104, 92) /bd:[ Ti0>A(26/104) Ti1>B(75/104) Li0>Cin(56/92) Bo0<S(53/104) Ro0<Cout(59/92) ]
input B;    //: /sn:0 {0}(373,159)(418,159){1}
//: {2}(422,159)(433,159)(433,141)(441,141){3}
//: {4}(420,161)(420,203){5}
//: {6}(422,205)(442,205){7}
//: {8}(420,207)(420,257)(442,257){9}
input A;    //: /sn:0 {0}(371,136)(410,136){1}
//: {2}(414,136)(441,136){3}
//: {4}(412,138)(412,198){5}
//: {6}(414,200)(442,200){7}
//: {8}(412,202)(412,225)(442,225){9}
input Cin;    //: /sn:0 {0}(371,177)(396,177){1}
//: {2}(400,177)(509,177)(509,156)(515,156){3}
//: {4}(398,179)(398,228){5}
//: {6}(400,230)(442,230){7}
//: {8}(398,232)(398,262)(442,262){9}
output Cout;    //: /sn:0 /dp:1 {0}(579,246)(617,246){1}
output S;    //: /sn:0 /dp:1 {0}(536,154)(597,154){1}
wire w13;    //: /sn:0 {0}(539,206)(548,206)(548,243)(558,243){1}
wire w3;    //: /sn:0 {0}(463,203)(518,203){1}
wire w12;    //: /sn:0 /dp:1 {0}(518,208)(473,208)(473,228)(463,228){1}
wire w2;    //: /sn:0 {0}(462,139)(505,139)(505,151)(515,151){1}
wire w15;    //: /sn:0 /dp:1 {0}(558,248)(473,248)(473,260)(463,260){1}
//: enddecls

  and g8 (.I0(B), .I1(Cin), .Z(w15));   //: @(453,260) /sn:0 /delay:" 2" /w:[ 9 9 1 ]
  xor g4 (.I0(w2), .I1(Cin), .Z(S));   //: @(526,154) /sn:0 /delay:" 3" /w:[ 1 3 0 ]
  //: joint g16 (Cin) @(398, 230) /w:[ 6 5 -1 8 ]
  xor g3 (.I0(A), .I1(B), .Z(w2));   //: @(452,139) /sn:0 /delay:" 3" /w:[ 3 3 0 ]
  //: output g17 (Cout) @(614,246) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(369,177) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(371,159) /sn:0 /w:[ 0 ]
  or g10 (.I0(w13), .I1(w15), .Z(Cout));   //: @(569,246) /sn:0 /delay:" 2" /w:[ 1 0 0 ]
  and g6 (.I0(A), .I1(B), .Z(w3));   //: @(453,203) /sn:0 /delay:" 2" /w:[ 7 7 0 ]
  or g9 (.I0(w3), .I1(w12), .Z(w13));   //: @(529,206) /sn:0 /delay:" 2" /w:[ 1 0 0 ]
  and g7 (.I0(A), .I1(Cin), .Z(w12));   //: @(453,228) /sn:0 /delay:" 2" /w:[ 9 7 1 ]
  //: joint g12 (B) @(420, 159) /w:[ 2 -1 1 4 ]
  //: joint g14 (Cin) @(398, 177) /w:[ 2 -1 1 4 ]
  //: joint g11 (A) @(412, 136) /w:[ 2 -1 1 4 ]
  //: output g5 (S) @(594,154) /sn:0 /w:[ 1 ]
  //: joint g15 (B) @(420, 205) /w:[ 6 5 -1 8 ]
  //: input g0 (A) @(369,136) /sn:0 /w:[ 0 ]
  //: joint g13 (A) @(412, 200) /w:[ 6 5 -1 8 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(166,174)(245,174){1}
wire w7;    //: /sn:0 {0}(342,60)(321,60)(321,117){1}
wire w4;    //: /sn:0 {0}(351,177)(391,177){1}
wire w5;    //: /sn:0 {0}(248,60)(272,60)(272,117){1}
wire w9;    //: /sn:0 {0}(299,249)(299,211){1}
//: enddecls

  led g4 (.I(w4));   //: @(398,177) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: switch g3 (w7) @(360,60) /sn:0 /R:2 /w:[ 0 ] /st:1
  //: switch g2 (w6) @(149,174) /sn:0 /w:[ 0 ] /st:1
  //: switch g1 (w5) @(231,60) /sn:0 /w:[ 0 ] /st:1
  led g5 (.I(w9));   //: @(299,256) /sn:0 /R:2 /w:[ 0 ] /type:0
  full_adder g0 (.B(w7), .A(w5), .Cin(w6), .S(w9), .Cout(w4));   //: @(246, 118) /sz:(104, 92) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<1 Ro0<0 ]

endmodule
