//: version "1.8.7"

module PFA(Cin, B, P, S, A, G);
//: interface  /sz:(52, 47) /bd:[ Ti0>A(9/52) Ti1>B(39/52) Ri0>Cin(24/47) Bo0<S(40/52) Bo1<P(7/52) Bo2<G(18/52) ]
input B;    //: /sn:0 /dp:1 {0}(214,137)(104,137){1}
//: {2}(102,135)(102,66){3}
//: {4}(104,64)(139,64){5}
//: {6}(100,64)(84,64)(84,80)(76,80){7}
//: {8}(102,139)(102,163)(212,163){9}
input A;    //: /sn:0 /dp:1 {0}(139,59)(129,59){1}
//: {2}(125,59)(76,59){3}
//: {4}(127,61)(127,130){5}
//: {6}(129,132)(214,132){7}
//: {8}(127,134)(127,158)(212,158){9}
output G;    //: /sn:0 {0}(283,161)(233,161){1}
input Cin;    //: /sn:0 {0}(76,104)(209,104)(209,74)(219,74){1}
output P;    //: /sn:0 {0}(283,135)(235,135){1}
output S;    //: /sn:0 /dp:1 {0}(240,72)(283,72){1}
wire w2;    //: /sn:0 {0}(160,62)(209,62)(209,69)(219,69){1}
//: enddecls

  xor g4 (.I0(w2), .I1(Cin), .Z(S));   //: @(230,72) /sn:0 /delay:" 3" /w:[ 1 1 0 ]
  //: joint g8 (A) @(127, 59) /w:[ 1 -1 2 4 ]
  xor g3 (.I0(A), .I1(B), .Z(w2));   //: @(150,62) /sn:0 /delay:" 3" /w:[ 0 5 0 ]
  //: input g2 (Cin) @(74,104) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(74,80) /sn:0 /w:[ 7 ]
  //: joint g10 (A) @(127, 132) /w:[ 6 5 -1 8 ]
  and g6 (.I0(A), .I1(B), .Z(G));   //: @(223,161) /sn:0 /delay:" 2" /w:[ 9 9 1 ]
  or g7 (.I0(A), .I1(B), .Z(P));   //: @(225,135) /sn:0 /delay:" 2" /w:[ 7 0 1 ]
  //: joint g9 (B) @(102, 64) /w:[ 4 -1 6 3 ]
  //: output g12 (P) @(280,135) /sn:0 /w:[ 0 ]
  //: output g5 (S) @(280,72) /sn:0 /w:[ 1 ]
  //: joint g11 (B) @(102, 137) /w:[ 1 2 -1 8 ]
  //: input g0 (A) @(74,59) /sn:0 /w:[ 3 ]
  //: output g13 (G) @(280,161) /sn:0 /w:[ 0 ]

endmodule

module Carrylookahead_logic(P2, C1, G2, G0, C3, P0, C4, GG, G1, P1, P3, PG, G3, C2, C0);
//: interface  /sz:(196, 57) /bd:[ Ti0>G0(184/196) Ti1>P0(174/196) Ti2>G1(132/196) Ti3>P1(120/196) Ti4>G3(38/196) Ti5>P3(22/196) Ti6>P2(76/196) Ti7>G2(88/196) Ri0>C0(36/57) To0<C1(160/196) To1<C2(108/196) To2<C3(65/196) Lo0<C4(33/57) Bo0<GG(135/196) Bo1<PG(105/196) ]
input G2;    //: /sn:0 {0}(475,310)(472,310)(472,341)(184,341){1}
//: {2}(180,341)(61,341){3}
//: {4}(182,343)(182,476){5}
//: {6}(184,478)(358,478){7}
//: {8}(182,480)(182,641)(338,641){9}
input C0;    //: /sn:0 /dp:1 {0}(65,91)(324,91){1}
//: {2}(328,91)(338,91){3}
//: {4}(326,93)(326,144){5}
//: {6}(328,146)(341,146){7}
//: {8}(326,148)(326,236){9}
//: {10}(328,238)(358,238){11}
//: {12}(326,240)(326,370)(360,370){13}
output GG;    //: /sn:0 /dp:1 {0}(473,578)(537,578){1}
input P1;    //: /sn:0 {0}(360,380)(244,380){1}
//: {2}(242,378)(242,285){3}
//: {4}(244,283)(357,283){5}
//: {6}(242,281)(242,250){7}
//: {8}(244,248)(358,248){9}
//: {10}(242,246)(242,181){11}
//: {12}(244,179)(273,179){13}
//: {14}(242,177)(242,158){15}
//: {16}(244,156)(341,156){17}
//: {18}(240,156)(63,156){19}
//: {20}(242,382)(242,415){21}
//: {22}(244,417)(359,417){23}
//: {24}(242,419)(242,527){25}
//: {26}(244,529)(339,529){27}
//: {28}(242,531)(242,569)(337,569){29}
output C3;    //: /sn:0 /dp:1 {0}(496,302)(631,302){1}
output PG;    //: /sn:0 /dp:1 {0}(360,531)(454,531){1}
input G0;    //: /sn:0 /dp:1 {0}(65,122)(264,122){1}
//: {2}(268,122)(424,122){3}
//: {4}(266,124)(266,172){5}
//: {6}(268,174)(273,174){7}
//: {8}(266,176)(266,276){9}
//: {10}(268,278)(357,278){11}
//: {12}(266,280)(266,410){13}
//: {14}(268,412)(359,412){15}
//: {16}(266,414)(266,564)(337,564){17}
output C4;    //: /sn:0 {0}(612,446)(516,446){1}
output C2;    //: /sn:0 {0}(637,185)(448,185){1}
input P3;    //: /sn:0 {0}(338,612)(198,612){1}
//: {2}(196,610)(196,581){3}
//: {4}(198,579)(337,579){5}
//: {6}(196,577)(196,541){7}
//: {8}(198,539)(339,539){9}
//: {10}(196,537)(196,485){11}
//: {12}(198,483)(358,483){13}
//: {14}(196,481)(196,458){15}
//: {16}(198,456)(358,456){17}
//: {18}(196,454)(196,429){19}
//: {20}(198,427)(359,427){21}
//: {22}(196,425)(196,392){23}
//: {24}(198,390)(360,390){25}
//: {26}(194,390)(57,390){27}
//: {28}(196,614)(196,636)(338,636){29}
input G1;    //: /sn:0 {0}(62,190)(213,190){1}
//: {2}(217,190)(427,190){3}
//: {4}(215,192)(215,314){5}
//: {6}(217,316)(357,316){7}
//: {8}(215,318)(215,444){9}
//: {10}(217,446)(358,446){11}
//: {12}(215,448)(215,602)(338,602){13}
input G3;    //: /sn:0 {0}(452,586)(391,586)(391,657)(133,657)(133,501){1}
//: {2}(135,499)(487,499)(487,456)(495,456){3}
//: {4}(131,499)(64,499){5}
output C1;    //: /sn:0 /dp:1 {0}(445,120)(640,120){1}
input P0;    //: /sn:0 /dp:1 {0}(65,113)(85,113)(85,96)(309,96){1}
//: {2}(313,96)(338,96){3}
//: {4}(311,98)(311,149){5}
//: {6}(313,151)(341,151){7}
//: {8}(311,153)(311,241){9}
//: {10}(313,243)(358,243){11}
//: {12}(311,245)(311,373){13}
//: {14}(313,375)(360,375){15}
//: {16}(311,377)(311,524)(339,524){17}
input P2;    //: /sn:0 {0}(337,574)(228,574){1}
//: {2}(226,572)(226,536){3}
//: {4}(228,534)(339,534){5}
//: {6}(226,532)(226,453){7}
//: {8}(228,451)(358,451){9}
//: {10}(226,449)(226,424){11}
//: {12}(228,422)(359,422){13}
//: {14}(226,420)(226,387){15}
//: {16}(228,385)(360,385){17}
//: {18}(226,383)(226,313){19}
//: {20}(228,311)(357,311){21}
//: {22}(226,309)(226,290){23}
//: {24}(228,288)(357,288){25}
//: {26}(226,286)(226,255){27}
//: {28}(228,253)(358,253){29}
//: {30}(224,253)(52,253){31}
//: {32}(226,576)(226,607)(338,607){33}
wire w6;    //: /sn:0 /dp:1 {0}(452,576)(369,576)(369,607)(359,607){1}
wire w16;    //: /sn:0 {0}(452,581)(379,581)(379,639)(359,639){1}
wire w7;    //: /sn:0 {0}(381,380)(485,380)(485,436)(495,436){1}
wire w4;    //: /sn:0 /dp:1 {0}(427,180)(417,180)(417,151)(362,151){1}
wire w3;    //: /sn:0 /dp:1 {0}(475,300)(388,300)(388,283)(378,283){1}
wire w0;    //: /sn:0 /dp:1 {0}(424,117)(402,117)(402,94)(359,94){1}
wire w18;    //: /sn:0 /dp:1 {0}(452,571)(358,571){1}
wire w1;    //: /sn:0 /dp:1 {0}(427,185)(319,185)(319,177)(294,177){1}
wire w8;    //: /sn:0 /dp:1 {0}(495,441)(459,441)(459,419)(380,419){1}
wire w14;    //: /sn:0 {0}(495,446)(389,446)(389,451)(379,451){1}
wire w2;    //: /sn:0 /dp:1 {0}(475,295)(445,295)(445,245)(379,245){1}
wire w15;    //: /sn:0 {0}(495,451)(408,451)(408,481)(379,481){1}
wire w9;    //: /sn:0 {0}(475,305)(388,305)(388,314)(378,314){1}
//: enddecls

  //: joint g44 (G1) @(215, 316) /w:[ 6 5 -1 8 ]
  and g8 (.I0(C0), .I1(P0), .I2(P1), .Z(w4));   //: @(352,151) /sn:0 /delay:" 2" /w:[ 7 7 17 1 ]
  and g4 (.I0(C0), .I1(P0), .Z(w0));   //: @(349,94) /sn:0 /delay:" 2" /w:[ 3 3 1 ]
  //: input g16 (P2) @(50,253) /sn:0 /w:[ 31 ]
  and g47 (.I0(G2), .I1(P3), .Z(w15));   //: @(369,481) /sn:0 /delay:" 2" /w:[ 7 13 1 ]
  //: output g3 (C1) @(637,120) /sn:0 /w:[ 1 ]
  and g26 (.I0(P2), .I1(G1), .Z(w9));   //: @(368,314) /sn:0 /delay:" 2" /w:[ 21 7 1 ]
  //: input g17 (G2) @(59,341) /sn:0 /w:[ 3 ]
  //: input g2 (G0) @(63,122) /sn:0 /w:[ 0 ]
  //: output g30 (C3) @(628,302) /sn:0 /w:[ 1 ]
  //: joint g23 (G0) @(266, 174) /w:[ 6 5 -1 8 ]
  //: joint g39 (G0) @(266, 278) /w:[ 10 9 -1 12 ]
  //: joint g24 (P1) @(242, 248) /w:[ 8 10 -1 7 ]
  //: input g1 (P0) @(63,113) /sn:0 /w:[ 0 ]
  or g29 (.I0(w2), .I1(w3), .I2(w9), .I3(G2), .Z(C3));   //: @(486,302) /sn:0 /delay:" 2" /w:[ 0 0 0 0 0 ]
  //: joint g60 (P1) @(242, 529) /w:[ 26 25 -1 28 ]
  //: output g51 (C4) @(609,446) /sn:0 /w:[ 0 ]
  and g18 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .Z(w2));   //: @(369,245) /sn:0 /delay:" 2" /w:[ 11 11 9 29 1 ]
  or g70 (.I0(w18), .I1(w6), .I2(w16), .I3(G3), .Z(GG));   //: @(463,578) /sn:0 /delay:" 2" /w:[ 0 0 0 0 0 ]
  //: joint g25 (P2) @(226, 253) /w:[ 28 -1 30 27 ]
  //: joint g10 (C0) @(326, 91) /w:[ 2 -1 1 4 ]
  //: joint g65 (P2) @(226, 574) /w:[ 1 2 -1 32 ]
  //: joint g64 (G1) @(215, 446) /w:[ 10 9 -1 12 ]
  //: joint g49 (P3) @(196, 456) /w:[ 16 18 -1 15 ]
  //: output g72 (GG) @(534,578) /sn:0 /w:[ 1 ]
  or g50 (.I0(w7), .I1(w8), .I2(w14), .I3(w15), .I4(G3), .Z(C4));   //: @(506,446) /sn:0 /delay:" 2" /w:[ 1 0 0 0 3 1 ]
  //: input g6 (G1) @(60,190) /sn:0 /w:[ 0 ]
  //: joint g35 (P0) @(311, 243) /w:[ 10 9 -1 12 ]
  //: joint g9 (P0) @(311, 96) /w:[ 2 -1 1 4 ]
  //: input g7 (P1) @(61,156) /sn:0 /w:[ 19 ]
  //: joint g56 (P0) @(311, 375) /w:[ 14 13 -1 16 ]
  and g58 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w18));   //: @(348,571) /sn:0 /delay:" 2" /w:[ 17 29 0 5 1 ]
  //: joint g68 (P3) @(196, 612) /w:[ 1 2 -1 28 ]
  //: input g31 (P3) @(55,390) /sn:0 /w:[ 27 ]
  and g22 (.I0(G0), .I1(P1), .I2(P2), .Z(w3));   //: @(368,283) /sn:0 /delay:" 2" /w:[ 11 5 25 1 ]
  //: joint g59 (G0) @(266, 412) /w:[ 14 13 -1 16 ]
  //: joint g71 (G3) @(133, 499) /w:[ 2 -1 4 1 ]
  and g67 (.I0(P3), .I1(G2), .Z(w16));   //: @(349,639) /sn:0 /delay:" 2" /w:[ 29 9 1 ]
  //: joint g45 (P2) @(226, 422) /w:[ 12 14 -1 11 ]
  //: joint g41 (P2) @(226, 385) /w:[ 16 18 -1 15 ]
  //: joint g36 (P1) @(242, 283) /w:[ 4 6 -1 3 ]
  and g33 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .I4(P3), .Z(w7));   //: @(371,380) /sn:0 /delay:" 2" /w:[ 13 15 0 17 25 0 ]
  //: joint g54 (P2) @(226, 451) /w:[ 8 10 -1 7 ]
  //: joint g42 (P3) @(196, 390) /w:[ 24 -1 26 23 ]
  //: joint g40 (P1) @(242, 380) /w:[ 1 2 -1 20 ]
  and g52 (.I0(P0), .I1(P1), .I2(P2), .I3(P3), .Z(PG));   //: @(350,531) /sn:0 /delay:" 2" /w:[ 17 27 5 9 0 ]
  //: joint g69 (G2) @(182, 478) /w:[ 6 5 -1 8 ]
  //: joint g66 (P3) @(196, 579) /w:[ 4 6 -1 3 ]
  //: joint g12 (G0) @(266, 122) /w:[ 2 -1 1 4 ]
  //: joint g46 (P3) @(196, 427) /w:[ 20 22 -1 19 ]
  //: joint g34 (C0) @(326, 238) /w:[ 10 9 -1 12 ]
  //: joint g28 (G1) @(215, 190) /w:[ 2 -1 1 4 ]
  //: output g57 (PG) @(451,531) /sn:0 /w:[ 1 ]
  or g14 (.I0(w4), .I1(w1), .I2(G1), .Z(C2));   //: @(438,185) /sn:0 /delay:" 2" /w:[ 0 0 3 1 ]
  and g11 (.I0(G0), .I1(P1), .Z(w1));   //: @(284,177) /sn:0 /delay:" 2" /w:[ 7 13 1 ]
  or g5 (.I0(w0), .I1(G0), .Z(C1));   //: @(435,120) /sn:0 /delay:" 2" /w:[ 0 3 0 ]
  //: joint g21 (P1) @(242, 179) /w:[ 12 14 -1 11 ]
  //: joint g19 (C0) @(326, 146) /w:[ 6 5 -1 8 ]
  //: joint g61 (P2) @(226, 534) /w:[ 4 6 -1 3 ]
  //: input g32 (G3) @(62,499) /sn:0 /w:[ 5 ]
  //: joint g20 (P0) @(311, 151) /w:[ 6 5 -1 8 ]
  and g63 (.I0(G1), .I1(P2), .I2(P3), .Z(w6));   //: @(349,607) /sn:0 /delay:" 2" /w:[ 13 33 0 1 ]
  and g43 (.I0(G1), .I1(P2), .I2(P3), .Z(w14));   //: @(369,451) /sn:0 /delay:" 2" /w:[ 11 9 17 1 ]
  and g38 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w8));   //: @(370,419) /sn:0 /delay:" 2" /w:[ 15 23 13 21 1 ]
  //: output g15 (C2) @(634,185) /sn:0 /w:[ 0 ]
  //: input g0 (C0) @(63,91) /sn:0 /w:[ 0 ]
  //: joint g48 (G2) @(182, 341) /w:[ 1 -1 2 4 ]
  //: joint g27 (P2) @(226, 288) /w:[ 24 26 -1 23 ]
  //: joint g37 (P2) @(226, 311) /w:[ 20 22 -1 19 ]
  //: joint g62 (P3) @(196, 539) /w:[ 8 10 -1 7 ]
  //: joint g55 (P1) @(242, 417) /w:[ 22 21 -1 24 ]
  //: joint g13 (P1) @(242, 156) /w:[ 16 -1 18 15 ]
  //: joint g53 (P3) @(196, 483) /w:[ 12 14 -1 11 ]

endmodule

module Lookahead_Carry_Unit(G12, G4, P4, C0, P0, C16, GG, P8, P12, PG, G8, C4, C8, C12, G0);
//: interface  /sz:(697, 107) /bd:[ Ti0>G0(612/697) Ti1>P0(590/697) Ti2>G4(420/697) Ti3>P4(395/697) Ti4>G8(242/697) Ti5>P8(217/697) Ti6>G12(48/697) Ti7>P12(21/697) Ri0>C0(61/107) To0<C4(524/697) To1<C8(348/697) To2<C12(154/697) Lo0<C16(70/107) Bo0<PG(350/697) Bo1<GG(405/697) ]
input P4;    //: /sn:0 {0}(886,457)(694,457){1}
//: {2}(692,455)(692,371){3}
//: {4}(694,369)(885,369){5}
//: {6}(692,367)(692,338){7}
//: {8}(694,336)(885,336){9}
//: {10}(692,334)(692,275){11}
//: {12}(694,273)(881,273){13}
//: {14}(692,271)(692,237){15}
//: {16}(694,235)(878,235){17}
//: {18}(690,235)(680,235)(680,235)(83,235){19}
//: {20}(692,459)(692,503){21}
//: {22}(694,505)(886,505){23}
//: {24}(692,507)(692,699){25}
//: {26}(694,701)(889,701){27}
//: {28}(692,703)(692,762)(888,762){29}
output C12;    //: /sn:0 /dp:1 {0}(1026,398)(1130,398){1}
output GG;    //: /sn:0 /dp:1 {0}(1025,804)(1144,804){1}
input C0;    //: /sn:0 {0}(878,225)(823,225){1}
//: {2}(821,223)(821,92){3}
//: {4}(823,90)(882,90)(882,107)(892,107){5}
//: {6}(819,90)(92,90){7}
//: {8}(821,227)(821,324){9}
//: {10}(823,326)(885,326){11}
//: {12}(821,328)(821,447)(886,447){13}
input P8;    //: /sn:0 {0}(888,767)(645,767){1}
//: {2}(643,765)(643,708){3}
//: {4}(645,706)(889,706){5}
//: {6}(643,704)(643,549){7}
//: {8}(645,547)(885,547){9}
//: {10}(643,545)(643,512){11}
//: {12}(645,510)(886,510){13}
//: {14}(643,508)(643,464){15}
//: {16}(645,462)(886,462){17}
//: {18}(643,460)(643,394){19}
//: {20}(645,392)(883,392){21}
//: {22}(643,390)(643,376){23}
//: {24}(645,374)(885,374){25}
//: {26}(643,372)(643,343){27}
//: {28}(645,341)(885,341){29}
//: {30}(641,341)(93,341){31}
//: {32}(643,769)(643,796)(887,796){33}
input G8;    //: /sn:0 {0}(87,406)(491,406){1}
//: {2}(495,406)(1005,406){3}
//: {4}(493,408)(493,581){5}
//: {6}(495,583)(885,583){7}
//: {8}(493,585)(493,827)(884,827){9}
output C16;    //: /sn:0 /dp:1 {0}(1024,514)(1146,514){1}
output PG;    //: /sn:0 {0}(1139,703)(910,703){1}
input G0;    //: /sn:0 /dp:1 {0}(881,278)(736,278){1}
//: {2}(734,276)(734,141){3}
//: {4}(736,139)(982,139){5}
//: {6}(732,139)(93,139){7}
//: {8}(734,280)(734,362){9}
//: {10}(736,364)(885,364){11}
//: {12}(734,366)(734,498){13}
//: {14}(736,500)(886,500){15}
//: {16}(734,502)(734,757)(888,757){17}
output C4;    //: /sn:0 {0}(1146,137)(1003,137){1}
input G4;    //: /sn:0 {0}(80,304)(568,304)(568,305)(578,305){1}
//: {2}(582,305)(998,305)(998,275)(1000,275){3}
//: {4}(580,307)(580,395){5}
//: {6}(582,397)(883,397){7}
//: {8}(580,399)(580,540){9}
//: {10}(582,542)(885,542){11}
//: {12}(580,544)(580,791)(887,791){13}
input P12;    //: /sn:0 {0}(887,801)(553,801){1}
//: {2}(551,799)(551,774){3}
//: {4}(553,772)(888,772){5}
//: {6}(551,770)(551,713){7}
//: {8}(553,711)(889,711){9}
//: {10}(551,709)(551,590){11}
//: {12}(553,588)(885,588){13}
//: {14}(551,586)(551,554){15}
//: {16}(553,552)(885,552){17}
//: {18}(551,550)(551,517){19}
//: {20}(553,515)(886,515){21}
//: {22}(551,513)(551,469){23}
//: {24}(553,467)(886,467){25}
//: {26}(549,467)(86,467){27}
//: {28}(551,803)(551,832)(884,832){29}
input P0;    //: /sn:0 {0}(93,119)(783,119){1}
//: {2}(787,119)(882,119)(882,112)(892,112){3}
//: {4}(785,121)(785,228){5}
//: {6}(787,230)(878,230){7}
//: {8}(785,232)(785,329){9}
//: {10}(787,331)(885,331){11}
//: {12}(785,333)(785,450){13}
//: {14}(787,452)(886,452){15}
//: {16}(785,454)(785,696)(889,696){17}
output C8;    //: /sn:0 {0}(1139,270)(1021,270){1}
input G12;    //: /sn:0 {0}(1004,812)(980,812)(980,842)(371,842)(371,639){1}
//: {2}(373,637)(985,637)(985,524)(1003,524){3}
//: {4}(369,637)(108,637){5}
wire w16;    //: /sn:0 {0}(1004,807)(915,807)(915,830)(905,830){1}
wire w7;    //: /sn:0 {0}(907,457)(993,457)(993,504)(1003,504){1}
wire w4;    //: /sn:0 /dp:1 {0}(1005,396)(982,396)(982,369)(906,369){1}
wire w0;    //: /sn:0 /dp:1 {0}(982,134)(924,134)(924,110)(913,110){1}
wire w3;    //: /sn:0 /dp:1 {0}(1005,391)(990,391)(990,333)(906,333){1}
wire w18;    //: /sn:0 /dp:1 {0}(1004,802)(918,802)(918,796)(908,796){1}
wire w10;    //: /sn:0 /dp:1 {0}(1003,509)(917,509)(917,507)(907,507){1}
wire w1;    //: /sn:0 /dp:1 {0}(1000,265)(956,265)(956,230)(899,230){1}
wire w8;    //: /sn:0 {0}(904,395)(970,395)(970,401)(1005,401){1}
wire w14;    //: /sn:0 {0}(1003,514)(916,514)(916,547)(906,547){1}
wire w2;    //: /sn:0 /dp:1 {0}(1000,270)(912,270)(912,276)(902,276){1}
wire w15;    //: /sn:0 {0}(1003,519)(950,519)(950,586)(906,586){1}
wire w9;    //: /sn:0 {0}(909,764)(994,764)(994,797)(1004,797){1}
//: enddecls

  //: input g8 (G12) @(106,637) /sn:0 /w:[ 5 ]
  //: joint g44 (G4) @(580, 397) /w:[ 6 5 -1 8 ]
  //: input g4 (G4) @(78,304) /sn:0 /w:[ 0 ]
  //: input g3 (P4) @(81,235) /sn:0 /w:[ 19 ]
  //: joint g16 (P4) @(692, 235) /w:[ 16 -1 18 15 ]
  //: joint g47 (G8) @(493, 406) /w:[ 2 -1 1 4 ]
  //: joint g17 (G0) @(734, 139) /w:[ 4 -1 6 3 ]
  //: joint g26 (G0) @(734, 278) /w:[ 1 2 -1 8 ]
  //: input g2 (C0) @(90,90) /sn:0 /w:[ 7 ]
  //: joint g23 (P4) @(692, 273) /w:[ 12 14 -1 11 ]
  //: joint g30 (P8) @(643, 374) /w:[ 24 26 -1 23 ]
  //: input g1 (P0) @(91,119) /sn:0 /w:[ 0 ]
  and g24 (.I0(G0), .I1(P4), .I2(P8), .Z(w4));   //: @(896,369) /sn:0 /delay:" 2" /w:[ 11 5 25 1 ]
  //: joint g39 (G0) @(734, 364) /w:[ 10 9 -1 12 ]
  //: joint g29 (C0) @(821, 326) /w:[ 10 9 -1 12 ]
  //: joint g60 (P4) @(692, 701) /w:[ 26 25 -1 28 ]
  //: output g51 (C16) @(1143,514) /sn:0 /w:[ 1 ]
  or g18 (.I0(w1), .I1(w2), .I2(G4), .Z(C8));   //: @(1011,270) /sn:0 /delay:" 2" /w:[ 0 0 3 1 ]
  or g70 (.I0(w9), .I1(w18), .I2(w16), .I3(G12), .Z(GG));   //: @(1015,804) /sn:0 /delay:" 2" /w:[ 1 0 0 0 0 ]
  or g10 (.I0(w0), .I1(G0), .Z(C4));   //: @(993,137) /sn:0 /delay:" 2" /w:[ 0 5 1 ]
  //: joint g25 (P4) @(692, 336) /w:[ 8 10 -1 7 ]
  //: joint g65 (P8) @(643, 767) /w:[ 1 2 -1 32 ]
  //: joint g64 (G4) @(580, 542) /w:[ 10 9 -1 12 ]
  //: output g72 (GG) @(1141,804) /sn:0 /w:[ 1 ]
  or g49 (.I0(w7), .I1(w10), .I2(w14), .I3(w15), .I4(G12), .Z(C16));   //: @(1014,514) /sn:0 /delay:" 2" /w:[ 1 0 0 0 3 0 ]
  //: input g6 (P8) @(91,341) /sn:0 /w:[ 31 ]
  //: joint g50 (P12) @(551, 552) /w:[ 16 18 -1 15 ]
  and g9 (.I0(C0), .I1(P0), .Z(w0));   //: @(903,110) /sn:0 /delay:" 2" /w:[ 5 3 1 ]
  //: input g7 (P12) @(84,467) /sn:0 /w:[ 27 ]
  //: joint g35 (G4) @(580, 305) /w:[ 2 -1 1 4 ]
  //: joint g56 (P12) @(551, 588) /w:[ 12 14 -1 11 ]
  and g58 (.I0(G0), .I1(P4), .I2(P8), .I3(P12), .Z(w9));   //: @(899,764) /sn:0 /delay:" 2" /w:[ 17 29 0 5 0 ]
  //: joint g68 (G8) @(493, 583) /w:[ 6 5 -1 8 ]
  //: joint g71 (G12) @(371, 637) /w:[ 2 -1 4 1 ]
  //: joint g22 (P0) @(785, 230) /w:[ 6 5 -1 8 ]
  or g31 (.I0(w3), .I1(w4), .I2(w8), .I3(G8), .Z(C12));   //: @(1016,398) /sn:0 /delay:" 2" /w:[ 0 0 1 3 0 ]
  //: joint g59 (G0) @(734, 500) /w:[ 14 13 -1 16 ]
  and g67 (.I0(G8), .I1(P12), .Z(w16));   //: @(895,830) /sn:0 /delay:" 2" /w:[ 9 29 1 ]
  and g33 (.I0(P8), .I1(G4), .Z(w8));   //: @(894,395) /sn:0 /delay:" 2" /w:[ 21 7 0 ]
  //: joint g36 (P4) @(692, 369) /w:[ 4 6 -1 3 ]
  //: joint g41 (P8) @(643, 462) /w:[ 16 18 -1 15 ]
  //: joint g45 (P8) @(643, 510) /w:[ 12 14 -1 11 ]
  //: joint g54 (P4) @(692, 505) /w:[ 22 21 -1 24 ]
  //: joint g40 (P4) @(692, 457) /w:[ 1 2 -1 20 ]
  //: joint g42 (P12) @(551, 467) /w:[ 24 -1 26 23 ]
  and g52 (.I0(P0), .I1(P4), .I2(P8), .I3(P12), .Z(PG));   //: @(900,703) /sn:0 /delay:" 2" /w:[ 17 27 5 9 1 ]
  //: joint g69 (P12) @(551, 801) /w:[ 1 2 -1 28 ]
  //: joint g66 (P12) @(551, 772) /w:[ 4 6 -1 3 ]
  and g12 (.I0(C0), .I1(P0), .I2(P4), .Z(w1));   //: @(889,230) /sn:0 /delay:" 2" /w:[ 0 7 17 1 ]
  and g28 (.I0(C0), .I1(P0), .I2(P4), .I3(P8), .I4(P12), .Z(w7));   //: @(897,457) /sn:0 /delay:" 2" /w:[ 13 15 0 17 25 0 ]
  //: joint g34 (P0) @(785, 331) /w:[ 10 9 -1 12 ]
  and g46 (.I0(G8), .I1(P12), .Z(w15));   //: @(896,586) /sn:0 /delay:" 2" /w:[ 7 13 1 ]
  //: output g57 (PG) @(1136,703) /sn:0 /w:[ 0 ]
  //: input g5 (G8) @(85,406) /sn:0 /w:[ 0 ]
  //: output g11 (C4) @(1143,137) /sn:0 /w:[ 0 ]
  //: joint g14 (P0) @(785, 119) /w:[ 2 -1 1 4 ]
  //: output g19 (C8) @(1136,270) /sn:0 /w:[ 0 ]
  //: joint g21 (C0) @(821, 225) /w:[ 1 2 -1 8 ]
  //: joint g61 (P8) @(643, 706) /w:[ 4 6 -1 3 ]
  and g20 (.I0(C0), .I1(P0), .I2(P4), .I3(P8), .Z(w3));   //: @(896,333) /sn:0 /delay:" 2" /w:[ 11 11 9 29 1 ]
  //: output g32 (C12) @(1127,398) /sn:0 /w:[ 1 ]
  and g63 (.I0(G4), .I1(P8), .I2(P12), .Z(w18));   //: @(898,796) /sn:0 /delay:" 2" /w:[ 13 33 0 1 ]
  //: input g0 (G0) @(91,139) /sn:0 /w:[ 7 ]
  and g15 (.I0(P4), .I1(G0), .Z(w2));   //: @(892,276) /sn:0 /delay:" 2" /w:[ 13 0 1 ]
  and g38 (.I0(G0), .I1(P4), .I2(P8), .I3(P12), .Z(w10));   //: @(897,507) /sn:0 /delay:" 2" /w:[ 15 23 13 21 1 ]
  and g43 (.I0(G4), .I1(P8), .I2(P12), .Z(w14));   //: @(896,547) /sn:0 /delay:" 2" /w:[ 11 9 17 1 ]
  //: joint g27 (P8) @(643, 341) /w:[ 28 -1 30 27 ]
  //: joint g48 (P12) @(551, 515) /w:[ 20 22 -1 19 ]
  //: joint g37 (P8) @(643, 392) /w:[ 20 22 -1 19 ]
  //: joint g62 (P12) @(551, 711) /w:[ 8 10 -1 7 ]
  //: joint g55 (P8) @(643, 547) /w:[ 8 10 -1 7 ]
  //: joint g13 (C0) @(821, 90) /w:[ 4 -1 6 3 ]
  //: joint g53 (P0) @(785, 452) /w:[ 14 13 -1 16 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(619,442)(619,493)(543,493){1}
wire [15:0] w7;    //: /sn:0 {0}(591,150)(591,258){1}
wire w4;    //: /sn:0 {0}(490,460)(589,460)(589,442){1}
wire [15:0] w0;    //: /sn:0 {0}(691,151)(691,258){1}
wire w1;    //: /sn:0 {0}(451,355)(511,355)(511,354)(572,354){1}
wire w2;    //: /sn:0 {0}(845,359)(770,359){1}
wire [15:0] w5;    //: /sn:0 {0}(675,555)(675,442){1}
//: enddecls

  led g4 (.I(w4));   //: @(483,460) /sn:0 /R:1 /w:[ 0 ] /type:0
  led g3 (.I(w1));   //: @(444,355) /sn:0 /R:1 /w:[ 0 ] /type:0
  //: dip g2 (w0) @(691,141) /sn:0 /w:[ 0 ] /st:65535
  //: dip g1 (w7) @(591,140) /sn:0 /w:[ 0 ] /st:65535
  led g6 (.I(w5));   //: @(675,562) /sn:0 /R:2 /w:[ 0 ] /type:3
  //: switch g7 (w2) @(863,359) /sn:0 /R:2 /w:[ 0 ] /st:0
  led g5 (.I(w6));   //: @(536,493) /sn:0 /R:1 /w:[ 1 ] /type:0
  CLA16bits g0 (.B(w0), .A(w7), .Cin(w2), .Cout(w1), .G(w6), .P(w4), .S(w5));   //: @(573, 259) /sz:(196, 182) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 Bo1<1 Bo2<1 ]

endmodule

module CLA16bits(P, A, G, Cout, B, Cin, S);
//: interface  /sz:(196, 182) /bd:[ Ti0>A[15:0](18/196) Ti1>B[15:0](118/196) Ri0>Cin(100/182) Lo0<Cout(95/182) Bo0<S[15:0](102/196) Bo1<P(16/196) Bo2<G(46/196) ]
input [15:0] B;    //: /sn:0 {0}(1125,70)(1125,190)(953,190){1}
//: {2}(952,190)(770,190){3}
//: {4}(769,190)(590,190){5}
//: {6}(589,190)(401,190){7}
//: {8}(400,190)(364,190){9}
input [15:0] A;    //: /sn:0 {0}(1088,73)(1088,159)(878,159){1}
//: {2}(877,159)(688,159){3}
//: {4}(687,159)(509,159){5}
//: {6}(508,159)(311,159){7}
//: {8}(310,159)(280,159){9}
output G;    //: /sn:0 {0}(692,663)(692,619)(693,619)(693,575){1}
input Cin;    //: /sn:0 /dp:1 {0}(988,293)(1044,293)(1044,355){1}
//: {2}(1046,357)(1113,357){3}
//: {4}(1044,359)(1044,528)(986,528){5}
output Cout;    //: /sn:0 {0}(132,537)(287,537){1}
output P;    //: /sn:0 {0}(638,575)(638,620)(637,620)(637,665){1}
output [15:0] S;    //: /sn:0 /dp:1 {0}(158,412)(37,412){1}
wire w16;    //: /sn:0 /dp:1 {0}(442,466)(442,301)(428,301){1}
wire [3:0] w6;    //: /sn:0 {0}(592,234)(592,213)(590,213)(590,194){1}
wire w13;    //: /sn:0 {0}(637,235)(637,292)(671,292){1}
wire [3:0] w7;    //: /sn:0 {0}(878,225)(878,163){1}
wire w25;    //: /sn:0 {0}(335,347)(335,406)(336,406)(336,466){1}
wire w4;    //: /sn:0 {0}(230,242)(230,299)(297,299){1}
wire [3:0] w22;    //: /sn:0 {0}(313,234)(313,171)(311,171)(311,163){1}
wire [3:0] w3;    //: /sn:0 {0}(508,234)(508,200)(509,200)(509,163){1}
wire [3:0] w0;    //: /sn:0 /dp:1 {0}(164,397)(974,397)(974,340){1}
wire w20;    //: /sn:0 {0}(504,345)(504,405)(505,405)(505,466){1}
wire w30;    //: /sn:0 /dp:1 {0}(683,466)(683,402)(682,402)(682,339){1}
wire [3:0] w29;    //: /sn:0 /dp:1 {0}(164,427)(413,427)(413,347){1}
wire w12;    //: /sn:0 /dp:1 {0}(708,466)(708,402)(707,402)(707,339){1}
wire w18;    //: /sn:0 {0}(834,222)(834,291)(863,291){1}
wire w23;    //: /sn:0 {0}(529,345)(529,405)(530,405)(530,466){1}
wire [3:0] w10;    //: /sn:0 {0}(686,229)(686,200)(688,200)(688,163){1}
wire [3:0] w21;    //: /sn:0 {0}(400,234)(400,202)(401,202)(401,194){1}
wire [3:0] w1;    //: /sn:0 /dp:1 {0}(164,407)(783,407)(783,339){1}
wire w32;    //: /sn:0 /dp:1 {0}(878,466)(878,403)(877,403)(877,340){1}
wire [3:0] w8;    //: /sn:0 {0}(961,225)(961,200)(953,200)(953,194){1}
wire w17;    //: /sn:0 {0}(466,247)(466,298)(493,298){1}
wire [3:0] w14;    //: /sn:0 {0}(770,229)(770,194){1}
wire w2;    //: /sn:0 /dp:1 {0}(812,466)(812,294)(797,294){1}
wire [3:0] w11;    //: /sn:0 /dp:1 {0}(164,417)(605,417)(605,345){1}
wire w5;    //: /sn:0 /dp:1 {0}(900,466)(900,403)(899,403)(899,340){1}
wire w9;    //: /sn:0 /dp:1 {0}(636,466)(636,300)(619,300){1}
wire w26;    //: /sn:0 {0}(308,347)(308,406)(309,406)(309,466){1}
//: enddecls

  //: output g8 (P) @(637,662) /sn:0 /R:3 /w:[ 1 ]
  Lookahead_Carry_Unit g4 (.P12(w26), .G12(w25), .P8(w20), .G8(w23), .P4(w30), .G4(w12), .P0(w32), .G0(w5), .C0(Cin), .C12(w16), .C8(w9), .C4(w2), .C16(Cout), .GG(G), .PG(P));   //: @(288, 467) /sz:(697, 107) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>5 To0<0 To1<0 To2<0 Lo0<1 Bo0<1 Bo1<0 ]
  CLA g3 (.A(w22), .B(w21), .Cin(w16), .Cout(w4), .S(w29), .P(w26), .G(w25));   //: @(298, 235) /sz:(129, 111) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<1 Bo1<0 Bo2<0 ]
  tran g16(.Z(w14), .I(B[7:4]));   //: @(770,188) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  tran g17(.Z(w10), .I(A[7:4]));   //: @(688,157) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  CLA g2 (.B(w8), .A(w7), .Cin(Cin), .Cout(w18), .G(w5), .P(w32), .S(w0));   //: @(864, 226) /sz:(123, 113) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Bo0<1 Bo1<1 Bo2<1 ]
  led g23 (.I(w17));   //: @(466,240) /sn:0 /w:[ 0 ] /type:0
  led g24 (.I(w13));   //: @(637,228) /sn:0 /w:[ 0 ] /type:0
  CLA g1 (.B(w14), .A(w10), .Cin(w2), .Cout(w13), .G(w12), .P(w30), .S(w1));   //: @(672, 230) /sz:(124, 108) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<1 Bo1<1 Bo2<1 ]
  tran g18(.Z(w6), .I(B[11:8]));   //: @(590,188) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  led g25 (.I(w18));   //: @(834,215) /sn:0 /w:[ 0 ] /type:0
  //: input g10 (A) @(1088,71) /sn:0 /R:3 /w:[ 0 ]
  //: joint g6 (Cin) @(1044, 357) /w:[ 2 1 -1 4 ]
  //: output g9 (G) @(692,660) /sn:0 /R:3 /w:[ 0 ]
  //: output g7 (Cout) @(135,537) /sn:0 /R:2 /w:[ 0 ]
  led g22 (.I(w4));   //: @(230,235) /sn:0 /w:[ 0 ] /type:0
  tran g12(.Z(w22), .I(A[15:12]));   //: @(311,157) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  //: input g11 (B) @(1125,68) /sn:0 /R:3 /w:[ 0 ]
  //: input g5 (Cin) @(1115,357) /sn:0 /R:2 /w:[ 3 ]
  tran g14(.Z(w7), .I(A[3:0]));   //: @(878,157) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g19(.Z(w3), .I(A[11:8]));   //: @(509,157) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  //: output g21 (S) @(40,412) /sn:0 /R:2 /w:[ 1 ]
  concat g20 (.I0(w0), .I1(w1), .I2(w11), .I3(w29), .Z(S));   //: @(159,412) /sn:0 /R:2 /w:[ 0 0 0 0 0 ] /dr:0
  tran g15(.Z(w8), .I(B[3:0]));   //: @(953,188) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  CLA g0 (.B(w6), .A(w3), .Cin(w9), .Cout(w17), .G(w23), .P(w20), .S(w11));   //: @(494, 235) /sz:(124, 109) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<0 Bo1<0 Bo2<1 ]
  tran g13(.Z(w21), .I(B[15:12]));   //: @(401,188) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1

endmodule

module CLA(Cout, B, A, S, G, P, Cin);
//: interface  /sz:(129, 111) /bd:[ Ti0>A[3:0](15/129) Ti1>B[3:0](102/129) Ri0>Cin(66/111) Lo0<Cout(64/111) Bo0<S[3:0](115/129) Bo1<P(10/129) Bo2<G(37/129) ]
input [3:0] B;    //: /sn:0 {0}(91,36)(91,52)(180,52){1}
//: {2}(181,52)(276,52){3}
//: {4}(277,52)(378,52){5}
//: {6}(379,52)(470,52){7}
//: {8}(471,52)(509,52){9}
input [3:0] A;    //: /sn:0 {0}(68,37)(68,63)(151,63){1}
//: {2}(152,63)(245,63){3}
//: {4}(246,63)(346,63){5}
//: {6}(347,63)(443,63){7}
//: {8}(444,63)(452,63){9}
output G;    //: /sn:0 {0}(365,317)(365,276){1}
input Cin;    //: /sn:0 {0}(427,254)(498,254)(498,152){1}
//: {2}(500,150)(574,150){3}
//: {4}(498,148)(498,127)(488,127){5}
output Cout;    //: /sn:0 /dp:1 {0}(229,251)(144,251){1}
output P;    //: /sn:0 {0}(335,276)(335,317){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(97,203)(34,203){1}
wire w16;    //: /sn:0 {0}(358,156)(358,206)(362,206)(362,217){1}
wire w13;    //: /sn:0 {0}(379,106)(379,56){1}
wire w25;    //: /sn:0 {0}(295,103)(295,64)(277,64)(277,56){1}
wire w36;    //: /sn:0 {0}(192,154)(192,218)(103,218){1}
wire w22;    //: /sn:0 {0}(453,151)(453,207)(414,207)(414,217){1}
wire w0;    //: /sn:0 {0}(318,217)(318,164)(274,164)(274,153){1}
wire w3;    //: /sn:0 {0}(268,217)(268,182)(170,182)(170,154){1}
wire w20;    //: /sn:0 {0}(444,101)(444,67){1}
wire w30;    //: /sn:0 {0}(296,153)(296,208)(103,208){1}
wire w18;    //: /sn:0 {0}(380,156)(380,198)(103,198){1}
wire w19;    //: /sn:0 {0}(474,101)(474,64)(471,64)(471,56){1}
wire w23;    //: /sn:0 {0}(442,151)(442,192)(404,192)(404,217){1}
wire w10;    //: /sn:0 {0}(338,217)(338,129)(309,129){1}
wire w24;    //: /sn:0 {0}(475,151)(475,188)(103,188){1}
wire w31;    //: /sn:0 {0}(191,105)(191,66)(181,66)(181,56){1}
wire w1;    //: /sn:0 {0}(306,217)(306,170)(263,170)(263,153){1}
wire w32;    //: /sn:0 {0}(161,105)(161,87)(152,87)(152,67){1}
wire w17;    //: /sn:0 {0}(347,156)(347,207)(350,207)(350,217){1}
wire w14;    //: /sn:0 {0}(349,106)(349,75)(347,75)(347,67){1}
wire w2;    //: /sn:0 {0}(252,217)(252,192)(159,192)(159,154){1}
wire w11;    //: /sn:0 {0}(390,217)(390,168)(404,168)(404,132)(393,132){1}
wire w26;    //: /sn:0 {0}(265,103)(265,75)(246,75)(246,67){1}
wire w9;    //: /sn:0 {0}(295,217)(295,177)(250,177)(250,130)(205,130){1}
//: enddecls

  tran g8(.Z(w19), .I(B[0]));   //: @(471,50) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  PFA g4 (.A(w32), .B(w31), .Cin(w9), .S(w36), .P(w2), .G(w3));   //: @(152, 106) /sz:(52, 47) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<1 Bo2<1 ]
  //: joint g16 (Cin) @(498, 150) /w:[ 2 4 -1 1 ]
  PFA g3 (.A(w26), .B(w25), .Cin(w10), .S(w30), .P(w1), .G(w0));   //: @(256, 104) /sz:(52, 48) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<1 Bo2<1 ]
  //: output g17 (Cout) @(147,251) /sn:0 /R:2 /w:[ 1 ]
  PFA g2 (.A(w20), .B(w19), .Cin(Cin), .S(w24), .P(w23), .G(w22));   //: @(435, 102) /sz:(52, 48) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>5 Bo0<0 Bo1<0 Bo2<0 ]
  PFA g1 (.A(w14), .B(w13), .Cin(w11), .S(w18), .P(w17), .G(w16));   //: @(340, 107) /sz:(52, 48) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<0 ]
  concat g18 (.I0(w24), .I1(w18), .I2(w30), .I3(w36), .Z(S));   //: @(98,203) /sn:0 /R:2 /w:[ 1 1 1 1 0 ] /dr:0
  tran g10(.Z(w14), .I(A[1]));   //: @(347,61) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g6 (B) @(91,34) /sn:0 /R:3 /w:[ 0 ]
  tran g9(.Z(w13), .I(B[1]));   //: @(379,50) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g7(.Z(w20), .I(A[0]));   //: @(444,61) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g12(.Z(w26), .I(A[2]));   //: @(246,61) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g14(.Z(w32), .I(A[3]));   //: @(152,61) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g11(.Z(w25), .I(B[2]));   //: @(277,50) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: input g5 (A) @(68,35) /sn:0 /R:3 /w:[ 0 ]
  //: output g19 (S) @(37,203) /sn:0 /R:2 /w:[ 1 ]
  //: output g21 (G) @(365,314) /sn:0 /R:3 /w:[ 0 ]
  //: output g20 (P) @(335,314) /sn:0 /R:3 /w:[ 1 ]
  //: input g15 (Cin) @(576,150) /sn:0 /R:2 /w:[ 3 ]
  Carrylookahead_logic g0 (.G0(w22), .P0(w23), .G1(w16), .P1(w17), .G3(w3), .P3(w2), .P2(w1), .G2(w0), .C0(Cin), .C1(w11), .C2(w10), .C3(w9), .C4(Cout), .GG(G), .PG(P));   //: @(230, 218) /sz:(196, 57) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Ti3>1 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>0 To0<0 To1<0 To2<0 Lo0<0 Bo0<1 Bo1<0 ]
  tran g13(.Z(w31), .I(B[3]));   //: @(181,50) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1

endmodule
