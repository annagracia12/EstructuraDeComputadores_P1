//: version "1.8.7"

module half_adder(CO, S, B, A);
//: interface  /sz:(101, 76) /bd:[ Ti0>A(28/101) Ti1>B(64/101) Lo0<CO(38/76) Bo0<S(47/101) ]
input B;    //: /sn:0 {0}(348,356)(369,356){1}
//: {2}(373,356)(442,356)(442,251)(450,251){3}
//: {4}(371,358)(371,369)(453,369){5}
input A;    //: /sn:0 {0}(336,246)(402,246){1}
//: {2}(406,246)(450,246){3}
//: {4}(404,248)(404,364)(453,364){5}
output CO;    //: /sn:0 /dp:1 {0}(474,366)(523,366){1}
output S;    //: /sn:0 /dp:1 {0}(471,248)(522,248){1}
//: enddecls

  and g4 (.I0(B), .I1(A), .Z(CO));   //: @(464,366) /sn:0 /delay:" 2" /w:[ 5 5 0 ]
  //: output g3 (CO) @(520,366) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(519,248) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(346,356) /sn:0 /w:[ 0 ]
  //: joint g6 (A) @(404, 246) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(371, 356) /w:[ 2 -1 1 4 ]
  xor g5 (.I0(B), .I1(A), .Z(S));   //: @(461,248) /sn:0 /delay:" 3" /w:[ 3 3 0 ]
  //: input g0 (A) @(334,246) /sn:0 /w:[ 0 ]

endmodule

module SUMADOR_CPA(Cout, S, Cin, B0, A0);
//: interface  /sz:(165, 127) /bd:[ Ti0>A0[3:0](26/188) Ti1>B0[3:0](131/188) Ri0>Cin(57/127) Lo0<Cout(65/139) Bo0<S[3:0](92/188) ]
input [3:0] A0;    //: /sn:0 /dp:9 {0}(899,235)(815,235){1}
//: {2}(814,235)(675,235){3}
//: {4}(674,235)(532,235){5}
//: {6}(531,235)(390,235){7}
//: {8}(389,235)(264,235)(264,178){9}
input Cin;    //: /sn:0 {0}(295,317)(373,317){1}
output Cout;    //: /sn:0 /dp:1 {0}(896,304)(924,304){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(883,437)(933,437){1}
input [3:0] B0;    //: /sn:0 {0}(285,177)(285,223)(443,223){1}
//: {2}(444,223)(581,223){3}
//: {4}(582,223)(722,223){5}
//: {6}(723,223)(867,223){7}
//: {8}(868,223)(910,223){9}
wire w16;    //: /sn:0 {0}(877,452)(839,452)(839,347){1}
wire w6;    //: /sn:0 {0}(675,278)(675,239){1}
wire B;    //: /sn:0 {0}(443,279)(443,235)(444,235)(444,227){1}
wire w0;    //: /sn:0 {0}(871,275)(871,235)(868,235)(868,227){1}
wire A;    //: /sn:0 {0}(391,279)(391,247)(390,247)(390,239){1}
wire w12;    //: /sn:0 {0}(877,432)(552,432)(552,351){1}
wire w19;    //: /sn:0 {0}(468,308)(504,308)(504,317)(514,317){1}
wire w10;    //: /sn:0 {0}(584,279)(584,235)(582,235)(582,227){1}
wire w1;    //: /sn:0 {0}(819,275)(819,247)(815,247)(815,239){1}
wire w8;    //: /sn:0 {0}(877,422)(411,422)(411,351){1}
wire w14;    //: /sn:0 {0}(609,308)(647,308)(647,316)(657,316){1}
wire w11;    //: /sn:0 {0}(532,279)(532,239){1}
wire w15;    //: /sn:0 {0}(877,442)(695,442)(695,350){1}
wire w5;    //: /sn:0 {0}(727,278)(727,235)(723,235)(723,227){1}
wire w9;    //: /sn:0 /dp:1 {0}(752,307)(779,307)(779,313)(801,313){1}
//: enddecls

  tran g8(.Z(w6), .I(A0[2]));   //: @(675,233) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  //: output g4 (Cout) @(921,304) /sn:0 /w:[ 1 ]
  concat g16 (.I0(w8), .I1(w12), .I2(w15), .I3(w16), .Z(S));   //: @(882,437) /sn:0 /w:[ 0 0 0 0 0 ] /dr:1
  full_Adder g3 (.A(A), .B(B), .Cin(Cin), .S(w8), .Cout(w19));   //: @(374, 280) /sz:(93, 70) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<0 ]
  //: output g17 (S) @(930,437) /sn:0 /w:[ 1 ]
  full_Adder g2 (.A(w11), .B(w10), .Cin(w19), .S(w12), .Cout(w14));   //: @(515, 280) /sz:(93, 70) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<0 ]
  full_Adder g1 (.A(w6), .B(w5), .Cin(w14), .S(w15), .Cout(w9));   //: @(658, 279) /sz:(93, 70) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<0 ]
  //: input g10 (Cin) @(293,317) /sn:0 /w:[ 0 ]
  tran g6(.Z(A), .I(A0[0]));   //: @(390,233) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  tran g9(.Z(w1), .I(A0[3]));   //: @(815,233) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g7(.Z(w11), .I(A0[1]));   //: @(532,233) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  tran g12(.Z(B), .I(B0[0]));   //: @(444,221) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g14(.Z(w5), .I(B0[2]));   //: @(723,221) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g11 (B0) @(285,175) /sn:0 /R:3 /w:[ 0 ]
  //: input g5 (A0) @(264,176) /sn:0 /R:3 /w:[ 9 ]
  tran g15(.Z(w0), .I(B0[3]));   //: @(868,221) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  full_Adder g0 (.A(w1), .B(w0), .Cin(w9), .S(w16), .Cout(Cout));   //: @(802, 276) /sz:(93, 70) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<0 ]
  tran g13(.Z(w10), .I(B0[1]));   //: @(582,221) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1

endmodule

module full_Adder(Cout, Cin, B, S, A);
//: interface  /sz:(93, 70) /bd:[ Ti0>B(69/93) Ti1>A(17/93) Li0>Cin(37/70) Bo0<S(37/93) Ro0<Cout(28/70) ]
input B;    //: /sn:0 {0}(143,68)(187,68){1}
input A;    //: /sn:0 {0}(155,116)(177,116)(177,104)(187,104){1}
input Cin;    //: /sn:0 {0}(142,196)(333,196)(333,121)(357,121){1}
output Cout;    //: /sn:0 /dp:1 {0}(522,234)(628,234){1}
output S;    //: /sn:0 /dp:1 {0}(435,102)(567,102)(567,99)(577,99){1}
wire w3;    //: /sn:0 {0}(265,85)(357,85){1}
wire w8;    //: /sn:0 /dp:1 {0}(501,231)(396,231)(396,150){1}
wire w2;    //: /sn:0 {0}(226,133)(226,236)(501,236){1}
//: enddecls

  or g4 (.I0(w8), .I1(w2), .Z(Cout));   //: @(512,234) /sn:0 /delay:" 2" /w:[ 0 1 0 ]
  //: output g3 (Cout) @(625,234) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(140,196) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(141,68) /sn:0 /w:[ 0 ]
  half_adder g6 (.B(w3), .A(Cin), .CO(w8), .S(S));   //: @(358, 49) /sz:(76, 101) /sn:0 /p:[ Li0>1 Li1>1 Bo0<1 Ro0<0 ]
  //: output g7 (S) @(574,99) /sn:0 /w:[ 1 ]
  half_adder g5 (.B(B), .A(A), .CO(w2), .S(w3));   //: @(188, 32) /sz:(76, 101) /sn:0 /p:[ Li0>1 Li1>1 Bo0<0 Ro0<0 ]
  //: input g0 (A) @(153,116) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire [3:0] w4;    //: /sn:0 /dp:1 {0}(418,118)(418,196)(475,196)(475,206){1}
wire w3;    //: /sn:0 /dp:1 {0}(619,264)(687,264){1}
wire w1;    //: /sn:0 {0}(348,266)(452,266){1}
wire [3:0] w2;    //: /sn:0 {0}(533,335)(533,390)(532,390)(532,446){1}
wire [3:0] w5;    //: /sn:0 /dp:1 {0}(567,206)(567,126)(666,126)(666,103){1}
//: enddecls

  //: switch g4 (w3) @(705,264) /sn:0 /R:2 /w:[ 1 ] /st:1
  led g3 (.I(w1));   //: @(341,266) /sn:0 /R:1 /w:[ 0 ] /type:0
  //: dip g2 (w5) @(666,93) /sn:0 /w:[ 1 ] /st:15
  //: dip g1 (w4) @(418,108) /sn:0 /w:[ 0 ] /st:15
  led g5 (.I(w2));   //: @(532,453) /sn:0 /R:2 /w:[ 1 ] /type:3
  SUMADOR_CPA g0 (.B0(w5), .A0(w4), .Cin(w3), .Cout(w1), .S(w2));   //: @(453, 207) /sz:(165, 127) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Bo0<0 ]

endmodule
