//: version "1.8.7"

module CPA(A, S, B, Cout, Cin);
//: interface  /sz:(113, 80) /bd:[ Ti0>B[3:0](93/113) Ti1>A[3:0](26/113) Li0>Cin(49/80) Bo0<S[3:0](57/113) Ro0<Cout(50/80) ]
input [3:0] B;    //: /sn:0 {0}(50,34)(137,34){1}
//: {2}(138,34)(317,34){3}
//: {4}(318,34)(495,34){5}
//: {6}(496,34)(679,34){7}
//: {8}(680,34)(727,34){9}
input [3:0] A;    //: /sn:0 {0}(59,19)(88,19){1}
//: {2}(89,19)(262,19){3}
//: {4}(263,19)(446,19){5}
//: {6}(447,19)(629,19){7}
//: {8}(630,19)(717,19){9}
input Cin;    //: /sn:0 {0}(27,135)(63,135){1}
output Cout;    //: /sn:0 {0}(769,147)(710,147){1}
output [3:0] S;    //: /sn:0 {0}(384,326)(332,326)(332,294){1}
wire w16;    //: /sn:0 {0}(631,87)(631,31)(630,31)(630,23){1}
wire w13;    //: /sn:0 {0}(117,172)(117,268)(317,268)(317,288){1}
wire w6;    //: /sn:0 {0}(262,81)(262,31)(263,31)(263,23){1}
wire w4;    //: /sn:0 {0}(528,144)(604,144){1}
wire w3;    //: /sn:0 {0}(476,178)(476,244)(337,244)(337,288){1}
wire w0;    //: /sn:0 {0}(498,84)(498,46)(496,46)(496,38){1}
wire w18;    //: /sn:0 {0}(658,181)(658,268)(347,268)(347,288){1}
wire w10;    //: /sn:0 {0}(139,78)(139,46)(138,46)(138,38){1}
wire w1;    //: /sn:0 {0}(449,84)(449,27)(447,27)(447,23){1}
wire w8;    //: /sn:0 {0}(293,175)(293,248)(327,248)(327,288){1}
wire w14;    //: /sn:0 {0}(169,138)(231,138){1}
wire w11;    //: /sn:0 {0}(90,78)(90,31)(89,31)(89,23){1}
wire w15;    //: /sn:0 {0}(680,87)(680,38){1}
wire w5;    //: /sn:0 {0}(318,81)(318,38){1}
wire w9;    //: /sn:0 {0}(353,141)(422,141){1}
//: enddecls

  tran g8(.Z(w16), .I(A[3]));   //: @(630,17) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: input g4 (A) @(57,19) /sn:0 /w:[ 0 ]
  concat g16 (.I0(w13), .I1(w8), .I2(w3), .I3(w18), .Z(S));   //: @(332,293) /sn:0 /R:3 /w:[ 1 1 1 1 1 ] /dr:0
  full_adder g3 (.A(w16), .B(w15), .Cin(w4), .S(w18), .Cout(Cout));   //: @(605, 88) /sz:(104, 92) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<1 ]
  //: output g17 (S) @(381,326) /sn:0 /w:[ 0 ]
  full_adder g2 (.A(w11), .B(w10), .Cin(Cin), .S(w13), .Cout(w14));   //: @(64, 79) /sz:(104, 92) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<0 ]
  full_adder g1 (.A(w6), .B(w5), .Cin(w14), .S(w8), .Cout(w9));   //: @(232, 82) /sz:(120, 92) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<0 ]
  tran g10(.Z(w10), .I(B[0]));   //: @(138,32) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g6(.Z(w6), .I(A[1]));   //: @(263,17) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: input g9 (B) @(48,34) /sn:0 /w:[ 0 ]
  tran g7(.Z(w1), .I(A[2]));   //: @(447,17) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g12(.Z(w0), .I(B[2]));   //: @(496,32) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: output g14 (Cout) @(766,147) /sn:0 /w:[ 0 ]
  tran g11(.Z(w5), .I(B[1]));   //: @(318,32) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g5(.Z(w11), .I(A[0]));   //: @(89,17) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: input g15 (Cin) @(25,135) /sn:0 /w:[ 0 ]
  full_adder g0 (.A(w1), .B(w0), .Cin(w9), .S(w3), .Cout(w4));   //: @(423, 85) /sz:(104, 92) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<0 Ro0<0 ]
  tran g13(.Z(w15), .I(B[3]));   //: @(680,32) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1

endmodule

module full_adder(Cout, Cin, B, S, A);
//: interface  /sz:(104, 92) /bd:[ Ti0>B(75/104) Ti1>A(26/104) Li0>Cin(56/92) Bo0<S(53/104) Ro0<Cout(59/92) ]
input B;    //: /sn:0 {0}(373,159)(418,159){1}
//: {2}(422,159)(433,159)(433,141)(441,141){3}
//: {4}(420,161)(420,203){5}
//: {6}(422,205)(442,205){7}
//: {8}(420,207)(420,257)(442,257){9}
input A;    //: /sn:0 {0}(371,136)(410,136){1}
//: {2}(414,136)(441,136){3}
//: {4}(412,138)(412,198){5}
//: {6}(414,200)(442,200){7}
//: {8}(412,202)(412,225)(442,225){9}
input Cin;    //: /sn:0 {0}(371,177)(396,177){1}
//: {2}(400,177)(509,177)(509,156)(515,156){3}
//: {4}(398,179)(398,228){5}
//: {6}(400,230)(442,230){7}
//: {8}(398,232)(398,262)(442,262){9}
output Cout;    //: /sn:0 /dp:1 {0}(579,246)(617,246){1}
output S;    //: /sn:0 /dp:1 {0}(536,154)(597,154){1}
wire w13;    //: /sn:0 {0}(539,206)(548,206)(548,243)(558,243){1}
wire w3;    //: /sn:0 {0}(463,203)(518,203){1}
wire w12;    //: /sn:0 /dp:1 {0}(518,208)(473,208)(473,228)(463,228){1}
wire w2;    //: /sn:0 {0}(462,139)(505,139)(505,151)(515,151){1}
wire w15;    //: /sn:0 /dp:1 {0}(558,248)(473,248)(473,260)(463,260){1}
//: enddecls

  xor g4 (.I0(w2), .I1(Cin), .Z(S));   //: @(526,154) /sn:0 /delay:" 3" /w:[ 1 3 0 ]
  and g8 (.I0(B), .I1(Cin), .Z(w15));   //: @(453,260) /sn:0 /delay:" 2" /w:[ 9 9 1 ]
  xor g3 (.I0(A), .I1(B), .Z(w2));   //: @(452,139) /sn:0 /delay:" 3" /w:[ 3 3 0 ]
  //: joint g16 (Cin) @(398, 230) /w:[ 6 5 -1 8 ]
  //: output g17 (Cout) @(614,246) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(369,177) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(371,159) /sn:0 /w:[ 0 ]
  or g10 (.I0(w13), .I1(w15), .Z(Cout));   //: @(569,246) /sn:0 /delay:" 2" /w:[ 1 0 0 ]
  and g6 (.I0(A), .I1(B), .Z(w3));   //: @(453,203) /sn:0 /delay:" 2" /w:[ 7 7 0 ]
  and g7 (.I0(A), .I1(Cin), .Z(w12));   //: @(453,228) /sn:0 /delay:" 2" /w:[ 9 7 1 ]
  or g9 (.I0(w3), .I1(w12), .Z(w13));   //: @(529,206) /sn:0 /delay:" 2" /w:[ 1 0 0 ]
  //: joint g12 (B) @(420, 159) /w:[ 2 -1 1 4 ]
  //: output g5 (S) @(594,154) /sn:0 /w:[ 1 ]
  //: joint g11 (A) @(412, 136) /w:[ 2 -1 1 4 ]
  //: joint g14 (Cin) @(398, 177) /w:[ 2 -1 1 4 ]
  //: input g0 (A) @(369,136) /sn:0 /w:[ 0 ]
  //: joint g15 (B) @(420, 205) /w:[ 6 5 -1 8 ]
  //: joint g13 (A) @(412, 200) /w:[ 6 5 -1 8 ]

endmodule

module main;    //: root_module
wire [3:0] w4;    //: /sn:0 {0}(772,379)(772,393)(771,393)(771,407){1}
wire w3;    //: /sn:0 {0}(665,346)(690,346)(690,347)(714,347){1}
wire [3:0] w1;    //: /sn:0 {0}(807,253)(807,275)(808,275)(808,297){1}
wire [3:0] w2;    //: /sn:0 {0}(689,255)(689,280)(741,280)(741,297){1}
wire w5;    //: /sn:0 {0}(861,347)(845,347)(845,348)(829,348){1}
//: enddecls

  //: dip g4 (w2) @(689,245) /sn:0 /w:[ 0 ] /st:15
  //: switch g3 (w3) @(648,346) /sn:0 /w:[ 0 ] /st:0
  led g2 (.I(w4));   //: @(771,414) /sn:0 /R:2 /w:[ 1 ] /type:3
  led g1 (.I(w5));   //: @(868,347) /sn:0 /R:3 /w:[ 0 ] /type:0
  //: dip g5 (w1) @(807,243) /sn:0 /w:[ 0 ] /st:0
  CPA g0 (.A(w2), .B(w1), .Cin(w3), .S(w4), .Cout(w5));   //: @(715, 298) /sz:(113, 80) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<1 ]

endmodule
