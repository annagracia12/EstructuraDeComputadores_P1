//: version "1.8.7"

module half_adder(CO, S, B, A);
//: interface  /sz:(101, 76) /bd:[ Ti0>B(64/101) Ti1>A(28/101) Lo0<CO(38/76) Bo0<S(47/101) ]
input B;    //: /sn:0 {0}(348,356)(369,356){1}
//: {2}(373,356)(442,356)(442,251)(450,251){3}
//: {4}(371,358)(371,369)(453,369){5}
input A;    //: /sn:0 {0}(336,246)(402,246){1}
//: {2}(406,246)(450,246){3}
//: {4}(404,248)(404,364)(453,364){5}
output CO;    //: /sn:0 /dp:1 {0}(474,366)(523,366){1}
output S;    //: /sn:0 /dp:1 {0}(471,248)(522,248){1}
//: enddecls

  and g4 (.I0(B), .I1(A), .Z(CO));   //: @(464,366) /sn:0 /delay:" 2" /w:[ 5 5 0 ]
  //: output g3 (CO) @(520,366) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(519,248) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(346,356) /sn:0 /w:[ 0 ]
  //: joint g6 (A) @(404, 246) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(371, 356) /w:[ 2 -1 1 4 ]
  xor g5 (.I0(B), .I1(A), .Z(S));   //: @(461,248) /sn:0 /delay:" 3" /w:[ 3 3 0 ]
  //: input g0 (A) @(334,246) /sn:0 /w:[ 0 ]

endmodule

module RCA(B, Z, A);
//: interface  /sz:(165, 142) /bd:[ Ti0>A[3:0](22/165) Ti1>B[3:0](131/165) Bo0<Z[7:0](76/165) ]
input [3:0] B;    //: /sn:0 {0}(1475,59)(1400,59){1}
//: {2}(1399,59)(1289,59){3}
//: {4}(1288,59)(1147,59){5}
//: {6}(1146,59)(1034,59){7}
//: {8}(1033,59)(950,59){9}
input [3:0] A;    //: /sn:0 /dp:9 {0}(893,140)(907,140){1}
//: {2}(908,140)(1066,140){3}
//: {4}(1067,140)(1247,140){5}
//: {6}(1248,140)(1354,140)(1354,140)(1384,140){7}
//: {8}(1385,140)(1488,140){9}
output [7:0] Z;    //: /sn:0 {0}(1599,882)(1471,882){1}
wire w6;    //: /sn:0 {0}(1067,144)(1067,150)(1070,150)(1070,202){1}
//: {2}(1068,204)(960,204)(960,278){3}
//: {4}(958,280)(875,280)(875,509){5}
//: {6}(873,511)(735,511)(735,727){7}
//: {8}(875,513)(875,524)(876,524)(876,535){9}
//: {10}(960,282)(960,294){11}
//: {12}(1070,206)(1070,221){13}
wire w13;    //: /sn:0 {0}(1289,63)(1289,69)(1291,69)(1291,188){1}
//: {2}(1289,190)(1126,190){3}
//: {4}(1122,190)(967,190){5}
//: {6}(963,190)(778,190)(778,298){7}
//: {8}(965,192)(965,294){9}
//: {10}(1124,192)(1124,243)(1125,243)(1125,294){11}
//: {12}(1291,192)(1291,295){13}
wire w16;    //: /sn:0 {0}(1074,391)(957,391)(957,390)(947,390){1}
wire w7;    //: /sn:0 {0}(1075,221)(1075,124){1}
//: {2}(1077,122)(1253,122){3}
//: {4}(1257,122)(1399,122){5}
//: {6}(1401,120)(1401,69)(1400,69)(1400,63){7}
//: {8}(1401,124)(1401,219){9}
//: {10}(1255,124)(1255,221){11}
//: {12}(1073,122)(913,122)(913,220){13}
wire w34;    //: /sn:0 {0}(879,556)(879,588)(814,588)(814,621){1}
wire w25;    //: /sn:0 {0}(1113,678)(1113,867)(1465,867){1}
wire w0;    //: /sn:0 {0}(1385,144)(1385,170)(1396,170)(1396,199){1}
//: {2}(1394,201)(1286,201)(1286,277){3}
//: {4}(1284,279)(1142,279)(1142,453){5}
//: {6}(1140,455)(1029,455)(1029,729){7}
//: {8}(1142,457)(1142,480)(1143,480)(1143,504){9}
//: {10}(1286,281)(1286,295){11}
//: {12}(1396,203)(1396,219){13}
wire w22;    //: /sn:0 {0}(776,319)(776,343)(772,343)(772,353){1}
wire w36;    //: /sn:0 {0}(681,663)(681,792)(688,792)(688,802){1}
wire w20;    //: /sn:0 {0}(963,315)(963,355)(933,355)(933,365){1}
wire w29;    //: /sn:0 {0}(937,648)(871,648)(871,646)(828,646){1}
wire w30;    //: /sn:0 /dp:1 {0}(957,673)(957,783)(963,783)(963,793){1}
wire w37;    //: /sn:0 {0}(671,555)(671,617){1}
wire w42;    //: /sn:0 {0}(788,828)(735,828)(735,827)(725,827){1}
wire w12;    //: /sn:0 {0}(1272,434)(1272,857)(1465,857){1}
wire w19;    //: /sn:0 {0}(1123,315)(1123,362)(1107,362)(1107,372){1}
wire w18;    //: /sn:0 {0}(1065,639)(1006,639)(1006,652)(984,652){1}
wire w10;    //: /sn:0 {0}(1224,395)(1121,395){1}
wire w23;    //: /sn:0 /dp:1 {0}(900,386)(853,386)(853,343)(808,343)(808,353){1}
wire w24;    //: /sn:0 {0}(920,411)(920,513)(947,513)(947,627){1}
wire w21;    //: /sn:0 {0}(791,431)(791,621){1}
wire w1;    //: /sn:0 {0}(1248,144)(1248,150)(1250,150)(1250,202){1}
//: {2}(1248,204)(1119,204)(1119,267){3}
//: {4}(1117,269)(1008,269)(1008,504){5}
//: {6}(1006,506)(901,506)(901,616)(880,616)(880,731){7}
//: {8}(1008,508)(1008,532){9}
//: {10}(1119,271)(1119,282)(1120,282)(1120,294){11}
//: {12}(1250,206)(1250,221){13}
wire w31;    //: /sn:0 {0}(801,667)(801,797)(798,797)(798,807){1}
wire w32;    //: /sn:0 {0}(1011,553)(1011,617)(970,617)(970,627){1}
wire w8;    //: /sn:0 {0}(1073,242)(1073,362)(1084,362)(1084,372){1}
wire w46;    //: /sn:0 /dp:1 {0}(698,848)(698,897)(1465,897){1}
wire w17;    //: /sn:0 /dp:1 {0}(1094,415)(1094,600){1}
wire w27;    //: /sn:0 {0}(781,642)(708,642){1}
wire w44;    //: /sn:0 {0}(678,823)(633,823)(633,827)(623,827){1}
wire w28;    //: /sn:0 {0}(1146,525)(1146,590)(1130,590)(1130,600){1}
wire w33;    //: /sn:0 {0}(1013,532)(1013,479){1}
//: {2}(1015,477)(1145,477){3}
//: {4}(1147,475)(1147,63){5}
//: {6}(1147,479)(1147,491)(1148,491)(1148,504){7}
//: {8}(1011,477)(882,477){9}
//: {10}(878,477)(673,477)(673,534){11}
//: {12}(880,479)(880,507)(881,507)(881,535){13}
wire w35;    //: /sn:0 {0}(661,638)(586,638)(586,802){1}
wire w14;    //: /sn:0 {0}(1289,316)(1289,356){1}
wire w45;    //: /sn:0 {0}(883,752)(883,801)(821,801)(821,807){1}
wire w49;    //: /sn:0 /dp:1 {0}(596,848)(596,907)(1465,907){1}
wire w2;    //: /sn:0 {0}(1399,240)(1399,847)(1465,847){1}
wire w11;    //: /sn:0 {0}(911,241)(911,355)(910,355)(910,365){1}
wire w41;    //: /sn:0 {0}(1032,750)(1032,784)(999,784)(999,793){1}
wire w48;    //: /sn:0 {0}(738,748)(738,775)(711,775)(711,802){1}
wire w47;    //: /sn:0 /dp:1 {0}(576,823)(566,823)(566,917)(1465,917){1}
wire w15;    //: /sn:0 {0}(743,392)(694,392)(694,617){1}
wire w5;    //: /sn:0 {0}(1253,242)(1253,356){1}
wire w38;    //: /sn:0 {0}(982,871)(982,877)(1465,877){1}
wire w43;    //: /sn:0 /dp:1 {0}(808,853)(808,887)(1465,887){1}
wire w9;    //: /sn:0 {0}(908,144)(908,204){1}
//: {2}(906,206)(773,206)(773,277){3}
//: {4}(771,279)(668,279)(668,502){5}
//: {6}(666,504)(606,504)(606,725){7}
//: {8}(668,506)(668,534){9}
//: {10}(773,281)(773,298){11}
//: {12}(908,208)(908,220){13}
wire w26;    //: /sn:0 {0}(934,832)(835,832){1}
wire w40;    //: /sn:0 /dp:1 {0}(1034,729)(1034,703){1}
//: {2}(1034,699)(1034,63){3}
//: {4}(1032,701)(887,701){5}
//: {6}(883,701)(742,701){7}
//: {8}(738,701)(611,701)(611,725){9}
//: {10}(740,703)(740,727){11}
//: {12}(885,703)(885,731){13}
wire w51;    //: /sn:0 {0}(609,746)(609,802){1}
//: enddecls

  //: joint g4 (w7) @(1401, 122) /w:[ -1 6 5 8 ]
  //: joint g8 (w7) @(1255, 122) /w:[ 4 -1 3 10 ]
  //: joint g44 (w33) @(880, 477) /w:[ 9 -1 10 12 ]
  half_adder g16 (.B(w14), .A(w5), .CO(w10), .S(w12));   //: @(1225, 357) /sz:(101, 76) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  tran g3(.Z(w7), .I(B[0]));   //: @(1400,57) /sn:0 /R:1 /w:[ 7 2 1 ] /ss:1
  and g47 (.I0(w0), .I1(w40), .Z(w41));   //: @(1032,740) /sn:0 /R:3 /delay:" 2" /w:[ 7 0 0 ]
  and g17 (.I0(w0), .I1(w13), .Z(w14));   //: @(1289,306) /sn:0 /R:3 /delay:" 2" /w:[ 11 13 0 ]
  //: joint g26 (w1) @(1250, 204) /w:[ -1 1 2 12 ]
  and g2 (.I0(w0), .I1(w7), .Z(w2));   //: @(1399,230) /sn:0 /R:3 /delay:" 2" /w:[ 13 9 0 ]
  //: joint g23 (w13) @(1124, 190) /w:[ 3 -1 4 10 ]
  //: joint g30 (w9) @(908, 206) /w:[ -1 1 2 12 ]
  //: input g1 (B) @(1477,59) /sn:0 /R:2 /w:[ 0 ]
  and g24 (.I0(w9), .I1(w13), .Z(w22));   //: @(776,309) /sn:0 /R:3 /delay:" 2" /w:[ 11 7 0 ]
  and g39 (.I0(w6), .I1(w33), .Z(w34));   //: @(879,546) /sn:0 /R:3 /delay:" 2" /w:[ 9 13 0 ]
  half_adder g29 (.B(w23), .A(w22), .CO(w15), .S(w21));   //: @(744, 354) /sz:(101, 76) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  //: joint g60 (w40) @(740, 701) /w:[ 7 -1 8 10 ]
  and g51 (.I0(w1), .I1(w40), .Z(w45));   //: @(883,742) /sn:0 /R:3 /delay:" 2" /w:[ 7 13 0 ]
  //: joint g18 (w0) @(1396, 201) /w:[ -1 1 2 12 ]
  tran g10(.Z(w13), .I(B[1]));   //: @(1289,57) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  //: joint g25 (w13) @(965, 190) /w:[ 5 -1 6 8 ]
  //: joint g49 (w0) @(1142, 455) /w:[ -1 5 6 8 ]
  and g6 (.I0(w6), .I1(w7), .Z(w8));   //: @(1073,232) /sn:0 /R:3 /delay:" 2" /w:[ 13 0 0 ]
  full_Adder g50 (.B(w45), .A(w31), .Cin(w26), .Cout(w42), .S(w43));   //: @(789, 808) /sz:(45, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  and g7 (.I0(w9), .I1(w7), .Z(w11));   //: @(911,231) /sn:0 /R:3 /delay:" 2" /w:[ 13 13 0 ]
  //: joint g9 (w7) @(1075, 122) /w:[ 2 -1 12 1 ]
  and g35 (.I0(w1), .I1(w33), .Z(w32));   //: @(1011,543) /sn:0 /R:3 /delay:" 2" /w:[ 9 0 0 ]
  //: joint g56 (w40) @(885, 701) /w:[ 5 -1 6 12 ]
  full_Adder g58 (.B(w51), .A(w35), .Cin(w44), .Cout(w47), .S(w49));   //: @(577, 803) /sz:(45, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  and g22 (.I0(w6), .I1(w13), .Z(w20));   //: @(963,305) /sn:0 /R:3 /delay:" 2" /w:[ 11 9 0 ]
  half_adder g31 (.B(w28), .A(w17), .CO(w18), .S(w25));   //: @(1066, 601) /sz:(101, 76) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  and g59 (.I0(w9), .I1(w40), .Z(w51));   //: @(609,736) /sn:0 /R:3 /delay:" 2" /w:[ 7 9 0 ]
  //: joint g33 (w0) @(1286, 279) /w:[ -1 3 4 10 ]
  //: joint g36 (w33) @(1147, 477) /w:[ -1 4 3 6 ]
  //: joint g41 (w6) @(960, 280) /w:[ -1 3 4 10 ]
  //: joint g45 (w9) @(773, 279) /w:[ -1 3 4 10 ]
  full_Adder g54 (.B(w48), .A(w36), .Cin(w42), .Cout(w44), .S(w46));   //: @(679, 803) /sz:(45, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g40 (w33) @(1013, 477) /w:[ 2 -1 8 1 ]
  full_Adder g42 (.B(w15), .A(w37), .Cin(w27), .Cout(w35), .S(w36));   //: @(662, 618) /sz:(45, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g52 (w40) @(1034, 701) /w:[ -1 2 4 1 ]
  tran g12(.Z(w0), .I(A[0]));   //: @(1385,138) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: joint g28 (w6) @(1070, 204) /w:[ -1 1 2 12 ]
  full_Adder g34 (.B(w32), .A(w24), .Cin(w18), .Cout(w29), .S(w30));   //: @(938, 628) /sz:(45, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  half_adder g46 (.B(w41), .A(w30), .CO(w26), .S(w38));   //: @(935, 794) /sz:(101, 76) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  //: joint g57 (w6) @(875, 511) /w:[ -1 5 6 8 ]
  and g5 (.I0(w1), .I1(w7), .Z(w5));   //: @(1253,232) /sn:0 /R:3 /delay:" 2" /w:[ 13 11 0 ]
  tran g14(.Z(w6), .I(A[2]));   //: @(1067,138) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g11(.Z(w33), .I(B[2]));   //: @(1147,57) /sn:0 /R:1 /w:[ 5 6 5 ] /ss:1
  full_Adder g19 (.B(w19), .A(w8), .Cin(w10), .Cout(w16), .S(w17));   //: @(1075, 373) /sz:(45, 41) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g21 (w13) @(1291, 190) /w:[ -1 1 2 12 ]
  //: joint g61 (w9) @(668, 504) /w:[ -1 5 6 8 ]
  and g20 (.I0(w1), .I1(w13), .Z(w19));   //: @(1123,305) /sn:0 /R:3 /delay:" 2" /w:[ 11 11 0 ]
  and g32 (.I0(w0), .I1(w33), .Z(w28));   //: @(1146,515) /sn:0 /R:3 /delay:" 2" /w:[ 9 7 0 ]
  //: output g63 (Z) @(1596,882) /sn:0 /w:[ 0 ]
  //: input g0 (A) @(1490,140) /sn:0 /R:2 /w:[ 9 ]
  tran g15(.Z(w9), .I(A[3]));   //: @(908,138) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  full_Adder g38 (.B(w34), .A(w21), .Cin(w29), .Cout(w27), .S(w31));   //: @(782, 622) /sz:(45, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  and g43 (.I0(w9), .I1(w33), .Z(w37));   //: @(671,545) /sn:0 /R:3 /delay:" 2" /w:[ 9 11 0 ]
  full_Adder g27 (.B(w20), .A(w11), .Cin(w16), .Cout(w23), .S(w24));   //: @(901, 366) /sz:(45, 44) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  tran g48(.Z(w40), .I(B[3]));   //: @(1034,57) /sn:0 /R:1 /w:[ 3 8 7 ] /ss:1
  //: joint g37 (w1) @(1119, 269) /w:[ -1 3 4 10 ]
  concat g62 (.I0(w2), .I1(w12), .I2(w25), .I3(w38), .I4(w43), .I5(w46), .I6(w49), .I7(w47), .Z(Z));   //: @(1470,882) /sn:0 /w:[ 1 1 1 1 1 1 1 1 1 ] /dr:1
  and g55 (.I0(w6), .I1(w40), .Z(w48));   //: @(738,738) /sn:0 /R:3 /delay:" 2" /w:[ 7 11 0 ]
  tran g13(.Z(w1), .I(A[1]));   //: @(1248,138) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: joint g53 (w1) @(1008, 506) /w:[ -1 5 6 8 ]

endmodule

module full_Adder(Cin, B, Cout, S, A);
//: interface  /sz:(45, 44) /bd:[ Ti0>B(32/45) Ti1>A(9/45) Ri0>Cin(24/44) Lo0<Cout(20/44) Bo0<S(19/45) ]
input B;    //: /sn:0 {0}(85,83)(157,83)(157,71)(167,71){1}
input A;    //: /sn:0 {0}(86,50)(167,50){1}
input Cin;    //: /sn:0 {0}(84,123)(295,123)(295,82)(305,82){1}
output Cout;    //: /sn:0 /dp:1 {0}(401,160)(442,160){1}
output S;    //: /sn:0 /dp:1 {0}(357,72)(437,72){1}
wire w4;    //: /sn:0 {0}(331,103)(331,157)(380,157){1}
wire w3;    //: /sn:0 {0}(223,61)(305,61){1}
wire w2;    //: /sn:0 {0}(195,92)(195,162)(380,162){1}
//: enddecls

  half_adder g4 (.B(Cin), .A(w3), .CO(w4), .S(S));   //: @(306, 46) /sz:(50, 57) /sn:0 /p:[ Li0>1 Li1>1 Bo0<0 Ro0<0 ]
  half_adder g3 (.B(B), .A(A), .CO(w2), .S(w3));   //: @(168, 35) /sz:(54, 57) /sn:0 /p:[ Li0>1 Li1>1 Bo0<0 Ro0<0 ]
  //: input g2 (Cin) @(82,123) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(83,83) /sn:0 /w:[ 0 ]
  or g6 (.I0(w4), .I1(w2), .Z(Cout));   //: @(391,160) /sn:0 /delay:" 2" /w:[ 1 1 0 ]
  //: output g7 (Cout) @(439,160) /sn:0 /w:[ 1 ]
  //: output g5 (S) @(434,72) /sn:0 /w:[ 1 ]
  //: input g0 (A) @(84,50) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire [3:0] w3;    //: /sn:0 /dp:1 {0}(487,178)(487,274)(661,274)(661,281){1}
wire [3:0] w0;    //: /sn:0 /dp:1 {0}(802,172)(770,172)(770,281){1}
wire [7:0] w1;    //: /sn:0 {0}(735,493)(715,493)(715,425){1}
//: enddecls

  led g3 (.I(w1));   //: @(742,493) /sn:0 /R:3 /w:[ 0 ] /type:3
  //: dip g2 (w0) @(840,172) /sn:0 /R:3 /w:[ 0 ] /st:15
  //: dip g1 (w3) @(487,168) /sn:0 /w:[ 0 ] /st:11
  RCA g0 (.B(w0), .A(w3), .Z(w1));   //: @(639, 282) /sz:(165, 142) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 ]

endmodule
