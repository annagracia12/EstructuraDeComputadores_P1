//: version "1.8.7"

module half_adder(CO, S, B, A);
//: interface  /sz:(101, 76) /bd:[ Ti0>B(64/101) Ti1>A(28/101) Lo0<CO(38/76) Bo0<S(47/101) ]
input B;    //: /sn:0 {0}(348,356)(369,356){1}
//: {2}(373,356)(442,356)(442,251)(450,251){3}
//: {4}(371,358)(371,369)(453,369){5}
input A;    //: /sn:0 {0}(336,246)(402,246){1}
//: {2}(406,246)(450,246){3}
//: {4}(404,248)(404,364)(453,364){5}
output CO;    //: /sn:0 /dp:1 {0}(474,366)(523,366){1}
output S;    //: /sn:0 /dp:1 {0}(471,248)(522,248){1}
//: enddecls

  and g4 (.I0(B), .I1(A), .Z(CO));   //: @(464,366) /sn:0 /delay:" 2" /w:[ 5 5 0 ]
  //: output g3 (CO) @(520,366) /sn:0 /w:[ 1 ]
  //: output g2 (S) @(519,248) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(346,356) /sn:0 /w:[ 0 ]
  //: joint g6 (A) @(404, 246) /w:[ 2 -1 1 4 ]
  //: joint g7 (B) @(371, 356) /w:[ 2 -1 1 4 ]
  xor g5 (.I0(B), .I1(A), .Z(S));   //: @(461,248) /sn:0 /delay:" 3" /w:[ 3 3 0 ]
  //: input g0 (A) @(334,246) /sn:0 /w:[ 0 ]

endmodule

module full_Adder(Cout, Cin, B, S, A);
//: interface  /sz:(93, 70) /bd:[ Ti0>A(17/93) Ti1>B(69/93) Li0>Cin(37/70) Bo0<S(37/93) Ro0<Cout(28/70) ]
input B;    //: /sn:0 {0}(143,68)(187,68){1}
input A;    //: /sn:0 {0}(155,116)(177,116)(177,104)(187,104){1}
input Cin;    //: /sn:0 {0}(142,196)(333,196)(333,121)(357,121){1}
output Cout;    //: /sn:0 /dp:1 {0}(522,234)(628,234){1}
output S;    //: /sn:0 /dp:1 {0}(435,102)(567,102)(567,99)(577,99){1}
wire w3;    //: /sn:0 {0}(265,85)(357,85){1}
wire w8;    //: /sn:0 /dp:1 {0}(501,231)(396,231)(396,150){1}
wire w2;    //: /sn:0 {0}(226,133)(226,236)(501,236){1}
//: enddecls

  or g4 (.I0(w8), .I1(w2), .Z(Cout));   //: @(512,234) /sn:0 /delay:" 2" /w:[ 0 1 0 ]
  //: output g3 (Cout) @(625,234) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(140,196) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(141,68) /sn:0 /w:[ 0 ]
  half_adder g6 (.B(w3), .A(Cin), .CO(w8), .S(S));   //: @(358, 49) /sz:(76, 101) /sn:0 /p:[ Li0>1 Li1>1 Bo0<1 Ro0<0 ]
  //: output g7 (S) @(574,99) /sn:0 /w:[ 1 ]
  half_adder g5 (.B(B), .A(A), .CO(w2), .S(w3));   //: @(188, 32) /sz:(76, 101) /sn:0 /p:[ Li0>1 Li1>1 Bo0<0 Ro0<0 ]
  //: input g0 (A) @(153,116) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(155,235)(265,235)(265,244)(273,244){1}
wire w1;    //: /sn:0 /dp:1 {0}(343,206)(343,132)(389,132){1}
wire w8;    //: /sn:0 {0}(311,278)(311,323)(316,323)(316,332){1}
wire w5;    //: /sn:0 {0}(211,137)(252,137)(252,131){1}
//: {2}(254,129)(291,129)(291,206){3}
//: {4}(250,129)(242,129){5}
wire w9;    //: /sn:0 {0}(368,235)(430,235)(430,242)(443,242){1}
//: enddecls

  led g4 (.I(w8));   //: @(316,339) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: switch g3 (w1) @(407,132) /sn:0 /R:2 /w:[ 1 ] /st:1
  //: switch g2 (w6) @(138,235) /sn:0 /w:[ 0 ] /st:0
  //: switch g1 (w5) @(194,137) /sn:0 /w:[ 0 ] /st:1
  //: joint g6 (w5) @(252, 129) /w:[ 2 -1 4 1 ]
  led g5 (.I(w9));   //: @(450,242) /sn:0 /R:3 /w:[ 1 ] /type:0
  full_Adder g0 (.B(w1), .A(w5), .Cin(w6), .S(w8), .Cout(w9));   //: @(274, 207) /sz:(93, 70) /sn:0 /p:[ Ti0>0 Ti1>3 Li0>1 Bo0<0 Ro0<0 ]

endmodule
